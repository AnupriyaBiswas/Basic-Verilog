module and_gate (
    input wire A,
    input wire B,
    output wire Y
);

    and (Y, A, B);

endmodule
